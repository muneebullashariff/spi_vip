

	//Testbench top connects the DUV and the verification environment components

	//declare module

	//import uvm_pkg amd user_defined pkg


	//clock generation


	//instantiate duv

	//instantiate physical interface


	/*within initial block set the virtual interface,
	calling set config causes configuration settings to be created
	and placed in internal table of the component*/



	/*The UVM testbench is activated when the run_test() method is called,
	 the global run_test() task should be specified inside an initial block*/

	
