

	//Define type definition,functions and global variables for reuse

	//import uvm_pkg using scope resolution

	//include uvm_macros.svh

	//include all the tb component files
