
	/*agent_top that is sub-environment container that may contain one or
	more agents*/

	//extend agent_top class from uvm_env
	
	
	/*register with factory so can use create uvm_method and override in
	future if necessary*/


	//declare handle for agents to be created



	/*new constructor method that creates new component/object with
	leaf_instance "string name" and handle to its parent class*/
       


	/*build_phase necessary to get the automatic configuration of fields
	registered in the component by calling super.build_phase(phase)*/



	//create the agents
	


	//in runphase print topology
