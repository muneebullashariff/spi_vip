



	/*Efficient,reusable mechanism to organize configuration,extedned from
	uvm_object*/

	
	/*register with factory so can use create uvm_method and override in
	future if necessary*/

	

	//declare variables whether the env analysis components are used

	
	//declare variables if various agents are used

	
	//variable to tell if virtual_sequencer is present


	/*declare dynamic array of handles for the sub-component master and slave
	config classes*/
       

	//declare any variable to keep track of the transactions


	/*new constructor method that creates new component/object with
	leaf_instance "string name"*/	
	
	
