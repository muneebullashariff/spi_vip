


	/*Efficient,reusable mechanism to organize configuration,extedned from
	uvm_object*/

	
	/*register with factory so can use create uvm_method and override in
	future if necessary*/


 
	//declare handle for virtual interface
	

	//declare if the agent is active or passive
       

	//declare any variable to keep track of the transactions


	/*new constructor method that creates new component/object with
	leaf_instance "string name"*/	
	
