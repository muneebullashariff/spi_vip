



	/*transaction class holds the data_items\data_members required to drive
	stimulus to duv and also holds methods(task and functions) that manipulate those data_members 
	like copy,compare,could include constraints to generate meaningful data,could add print methods
	to print the data_members of the transaction class,extended from uvm_transaction or 
	uvm_sequence_item*/


	//declare class name extended from uvm_sequence_item
	
       
	/*register with factory so can use create uvm_method and override in
	future if necessary*/


	/*new constructor method that creates new component/object with
	leaf_instance "string name" and handle to its parent class*/


	/*constraints can be added to generate meaningful values according to
	the protocol*/


       //print method can be added to display the data_member values

