	
	/*A virtual sequence is a container to start multiple sequences
	on different sequencers in the environment*/

	/*extend virtual class from uvm_sequence parameterized with 
	uvm_sequence_item*/

	/*declare dynamic array of handle for master and slave
	sequencer*/

	//declare handle for virtual_sequencer

	//declare handle of all the sequences

	//declare handle for environment configuration class


	/*new constructor method that creates new component/object with
	leaf_instance "string name" and handle to its parent class*/

	

	/*build_phase necessary to get the automatic configuration of fields
	registered in the component by calling super.build_phase(phase)*/



	/*call get_config method,if value and the straing matches it returns
	the settings made with previous set call,if falied stop the simulation*/ 


	//initialize the dynamic arrays for master and slave sequencers


	/*assign master and slave sequencer handles tp virtual sequencer
	master and slave sequencer*/


	
