
	/*A virtual sequencer is used in the stimulus generation process
	to allow single sequences to control activity via several agents*/


	
	//declare dynamic array of handles for master and slave sequencer


	//declare handles for environment config class


	
	/*new constructor method that creates new component/object with
	leaf_instance "string name" and handle to its parent class*/

	

	/*build_phase necessary to get the automatic configuration of fields
	registered in the component by calling super.build_phase(phase)*/




	/*call get_config method,if value and the straing matches it returns
	the settings made with previous set call,if falied stop the simulation*/ 



	//create dynamic handles for master and slave sequencers	
