



	/*The sequencer control the flow of request and response sequence items between 
	sequences and the driver.Sequencer and driver uses TLM Interface to communicate transactions*/

	
	/*register with factory so can use create uvm_method and override in
	future if necessary*/


	/*new constructor method that creates new component/object with
	leaf_instance "string name"*/	
	
	
	
